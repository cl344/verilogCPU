module register0(out);
	output [31:0] out;
	out = 32'b0;
endmodule
