module andop(in1,in2,out);

input[31:0] in1,in2;
output[31:0] out;

and a0 (out[0 ],in1[0 ],in2[0 ]);
and a1 (out[1 ],in1[1 ],in2[1 ]);
and a2 (out[2 ],in1[2 ],in2[2 ]);
and a3 (out[3 ],in1[3 ],in2[3 ]);
and a4 (out[4 ],in1[4 ],in2[4 ]);
and a5 (out[5 ],in1[5 ],in2[5 ]);
and a6 (out[6 ],in1[6 ],in2[6 ]);
and a7 (out[7 ],in1[7 ],in2[7 ]);
and a8 (out[8 ],in1[8 ],in2[8 ]);
and a9 (out[9 ],in1[9 ],in2[9 ]);
and a10(out[10],in1[10],in2[10]);
and a11(out[11],in1[11],in2[11]);
and a12(out[12],in1[12],in2[12]);
and a13(out[13],in1[13],in2[13]);
and a14(out[14],in1[14],in2[14]);
and a15(out[15],in1[15],in2[15]);
and a16(out[16],in1[16],in2[16]);
and a17(out[17],in1[17],in2[17]);
and a18(out[18],in1[18],in2[18]);
and a19(out[19],in1[19],in2[19]);
and a20(out[20],in1[20],in2[20]);
and a21(out[21],in1[21],in2[21]);
and a22(out[22],in1[22],in2[22]);
and a23(out[23],in1[23],in2[23]);
and a24(out[24],in1[24],in2[24]);
and a25(out[25],in1[25],in2[25]);
and a26(out[26],in1[26],in2[26]);
and a27(out[27],in1[27],in2[27]);
and a28(out[28],in1[28],in2[28]);
and a29(out[29],in1[29],in2[29]);
and a30(out[30],in1[30],in2[30]);
and a31(out[31],in1[31],in2[31]);

endmodule
